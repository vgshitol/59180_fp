`timescale 1ns / 1ps

module Testbench;

	parameter CLOCK_PERIOD = 20;
	parameter MSG_LEN = 1024;
	//parameter MSG_LEN = 19;
	
	// INPUT REGISTERS
	reg clk; 
	reg resetn; 
	reg start;
	reg [7:0] msg;
	reg [11:0] msg_len; 

	// OUTPUT REGISTERS
	wire [7:0] hash;
	wire [7:0] hash_len; 
	wire valid;
	wire busy;

	// TB REGISTERS
	reg [8191:0] msg_str;
	reg [255:0] exp_hash_str;
	reg [255:0] obs_hash_str;
	reg cmp;

	reg  [255:0] test_vector [0:39] = {
		256'hEA152F2B47BCE24EFB66C479D4ADF17BD324D806E85FF75EE369EE50DC8F8BD1,
		256'h27921F8DDF392894460B70B3ED6C091E6421B7D2147DCD6031D7EFEBAD3030CC,
		256'hDD3F12E89DB41C61D3C05779705FA946A8C69C79EEFDC1B4A966A5F1AB35073D,
		256'h72ABD350DC287E8C4B95DD37BD796D79F90026C1BD4E0D99D2117BAAB26BC2CA,
		256'hA13AE46F62E433CE4CAD9E4F24C46F37B6B3815C8539A3659DAAECAAE1AB8FDB,
		256'h042383068C131A0D365B781DFCB20E855F4A68DE2072AA8D1E16181563D6F622,
		256'h415D3A751952454C1BB900700A2EB8C2814F0A30C34BC25CC37D3DE96159F4AE,
		256'h072F0834CC8FE7996E90ADED60228C18791E3A3DA38A3831DA880EDF7869909C,
		256'hC826D28C7F5BF948FBA9BB5EA028B4E377F1DE86EC5A2A1511BA4D692968EFD5,
		256'hD926F7E44B263CBA8F98E2A52B7BE175D406A2E81B462408BDBC408784C4284F,
		256'h98D44061E4D0EED4519061B947FD486B620F9B11CC3F4DF3F219E11E73B04FAD,
		256'hC23BF64CB9CE397460C685DE83EB40FE1B889CCDFDA5BE5DEA045AFCE30BB065,
		256'h4E55B9BA281BB67A05817083C3BFA219017E5DC455FD86C923641C922FFD67F2,
		256'h36CBE0424074FB55B2965FDE9FC305C88D142E97D82AC4B00974F68434733814,
		256'hD0FA0C36D76F9335615CE15E4A8B78C71B31F03DEA5EAB786CA91A887DA85DE4,
		256'hDB4C9CFE9D385D8CA329E27AEB495A0816C1AB051A57C231A134082661D71BED,
		256'h9EA695347CDDDFF9BC63ECE30FE231441D581768FE223DD6BD7367094FD216B3,
		256'h20593B39BB6D595019331601244411323F713085BB1A30218C972B96D9B7B7B3,
		256'h78C3560473F04C5DDE567433F1E125F417DD18518047D8D6B7B268620E78C19D,
		256'h9D8537BBA14AB9A9980CB4928274E6EBFDD7CBA1DAAE92F0750FD5B824B01362,
		256'h9BEBE7579EC1D075B6768AE981C54C7D60DB82931B074A618B0A68F84CBCCFE6,
		256'hD5B477858D82412D807BFBB60E6D770AF94D7B5537DEE497164673ED5C1A6D4F,
		256'h7562E4CF02443E85329C5ECE1294DF1DB8B52D44D052769C5F68987B0D7FC979,
		256'h511AD3AA185ACC22EB141A81C1EBDA05EADA4E0C07BFBAD3A4855DB3E96C2164,
		256'hE93B3C701C63199390D1D879AA68BA62D6677E03617B778C157D5FA2DFA382E8,
		256'h414825DCE3C8CE7CA480F15EB9BD765F10ECDB73EBC7C663967DA70B4E2A79F7,
		256'h5788DFE3C41A16A4CB06FC3C4E4BA39ADFFA3D1EEF04582E16A761B78BED1680,
		256'hAB5F4CB61A9F7C11600228695B771739CD00BC206B5CCA7FECD73B1C6B1B6781,
		256'h3529CCBE1165B6DF3EFF43B243207649D625017B897943846B1B95FDCCD8D300,
		256'hE300A2AF4B17DF61E1320BE0670177D4CE242A642047BB003FB50D8112497185,
		256'h5E8CBD381C53E6E26733255AAE669BBA2E42473E2D77064515C399D5AAEACB17,
		256'hB91E0C762169748D4E2B8D4972B63A4866CAAD1B5EBFB7F37DEADEB4424DF768,
		256'hCEBE4AFF9EAC2218017DDA5F8207BA830E989187256539BD7D31AE5E94FF0C6E,
		256'h249CFCCD50D66E722E80E79002CE3B302B4CA067483AB9CDEB474DBF555B7633,
		256'hA0AEF3C2B7AD6C45A3DE15D71767C7B432971532306454839F8BFF6E0DF5B97D,
		256'hB08F8899FEF00B282FDB550A4631A7989C568BAC2789480C8194522A17F01777,
		256'hF11AD59EE42A3969ADFAF398808FD1A2EFD1B4EDF686BE659A3DAB51F3839E83,
		256'h67D09BD54D5F9591CAA2535B1406E5B601D5F37C87BEA00EA86C2CF5385DA901,
		256'h8D55FABAB71392CE6A29B3A4FE185765AA7E5F2A829805CC306EE64CAFE3D25E,
		256'hD6C825A1BE1BCD24A2DCF1130D646BADE2C21CF6D48F043DCD46C01B80043FC1
	};
	
	//generate clock
	always #(CLOCK_PERIOD/2) clk = ~clk;

	// Instantiate the Unit Under Test (UUT)
	TOP dut (.clk(clk),.resetn(resetn),.start(start), .msg(msg), .msg_len(msg_len), 
		.hash(hash), .hash_len(hash_len), .valid(valid), .busy(busy));
	
	integer i=0,j=0,k=0;
	integer file,r;
		
	// Drive the testbench
	initial begin
		resetn=1'b1;
		clk = 1'b0;
		msg_str = 8192'h000102030405060708090A0B0C0D0E0F101112131415161718191A1B1C1D1E1F202122232425262728292A2B2C2D2E2F303132333435363738393A3B3C3D3E3F404142434445464748494A4B4C4D4E4F505152535455565758595A5B5C5D5E5F606162636465666768696A6B6C6D6E6F707172737475767778797A7B7C7D7E7F808182838485868788898A8B8C8D8E8F909192939495969798999A9B9C9D9E9FA0A1A2A3A4A5A6A7A8A9AAABACADAEAFB0B1B2B3B4B5B6B7B8B9BABBBCBDBEBFC0C1C2C3C4C5C6C7C8C9CACBCCCDCECFD0D1D2D3D4D5D6D7D8D9DADBDCDDDEDFE0E1E2E3E4E5E6E7E8E9EAEBECEDEEEFF0F1F2F3F4F5F6F7F8F9FAFBFCFDFEFF000102030405060708090A0B0C0D0E0F101112131415161718191A1B1C1D1E1F202122232425262728292A2B2C2D2E2F303132333435363738393A3B3C3D3E3F404142434445464748494A4B4C4D4E4F505152535455565758595A5B5C5D5E5F606162636465666768696A6B6C6D6E6F707172737475767778797A7B7C7D7E7F808182838485868788898A8B8C8D8E8F909192939495969798999A9B9C9D9E9FA0A1A2A3A4A5A6A7A8A9AAABACADAEAFB0B1B2B3B4B5B6B7B8B9BABBBCBDBEBFC0C1C2C3C4C5C6C7C8C9CACBCCCDCECFD0D1D2D3D4D5D6D7D8D9DADBDCDDDEDFE0E1E2E3E4E5E6E7E8E9EAEBECEDEEEFF0F1F2F3F4F5F6F7F8F9FAFBFCFDFEFF000102030405060708090A0B0C0D0E0F101112131415161718191A1B1C1D1E1F202122232425262728292A2B2C2D2E2F303132333435363738393A3B3C3D3E3F404142434445464748494A4B4C4D4E4F505152535455565758595A5B5C5D5E5F606162636465666768696A6B6C6D6E6F707172737475767778797A7B7C7D7E7F808182838485868788898A8B8C8D8E8F909192939495969798999A9B9C9D9E9FA0A1A2A3A4A5A6A7A8A9AAABACADAEAFB0B1B2B3B4B5B6B7B8B9BABBBCBDBEBFC0C1C2C3C4C5C6C7C8C9CACBCCCDCECFD0D1D2D3D4D5D6D7D8D9DADBDCDDDEDFE0E1E2E3E4E5E6E7E8E9EAEBECEDEEEFF0F1F2F3F4F5F6F7F8F9FAFBFCFDFEFF000102030405060708090A0B0C0D0E0F101112131415161718191A1B1C1D1E1F202122232425262728292A2B2C2D2E2F303132333435363738393A3B3C3D3E3F404142434445464748494A4B4C4D4E4F505152535455565758595A5B5C5D5E5F606162636465666768696A6B6C6D6E6F707172737475767778797A7B7C7D7E7F808182838485868788898A8B8C8D8E8F909192939495969798999A9B9C9D9E9FA0A1A2A3A4A5A6A7A8A9AAABACADAEAFB0B1B2B3B4B5B6B7B8B9BABBBCBDBEBFC0C1C2C3C4C5C6C7C8C9CACBCCCDCECFD0D1D2D3D4D5D6D7D8D9DADBDCDDDEDFE0E1E2E3E4E5E6E7E8E9EAEBECEDEEEFF0F1F2F3F4F5F6F7F8F9FAFBFCFDFEFF;
	    exp_hash_str = 256'hfcc4d63932d98c30cab597e60b7cca475bd9fbf984838c5cb5615c949f814615;
	   // msg_str = 8192'h000102030405060708090A0B0C0D0E0F101112;
	 	
	 	#(10*(CLOCK_PERIOD));
		resetn=1'b0;
		#(2*(CLOCK_PERIOD));
		
		resetn=1'b1;
		
		#(10*(CLOCK_PERIOD));
		for (j = 0; j < 40; j++) begin
			/* code */
			msg_len = j;
			exp_hash_str = test_vector[j];
		
			if(j==0) i = 0;
			else i = 1;

			#(5*CLOCK_PERIOD);
			start = 1;
			#(CLOCK_PERIOD);
			start = 0;

			while(i <=j ) begin
				load_msg();
			end 
			
			repeat(300) begin
				#((CLOCK_PERIOD));
			end	

		end

		$stop;
		
	end

	task load_msg;
    begin
	      if(~busy) begin 
	      	msg  = msg_str>>(1024-i)*8;
	      	i = i + 1;
	      end
	      else begin
	      	msg = msg;
	      	i = i;
	      end
	      #((CLOCK_PERIOD));
    end
  	endtask

	// Get the output string
	always@(posedge clk) begin
		if(~resetn) obs_hash_str <= 0;
		else if(valid==1'b1) begin
		//	 $display("VALID HIGH!");
			 obs_hash_str <= {obs_hash_str[247:0],hash};
		end
		else if(obs_hash_str==exp_hash_str) obs_hash_str <= 0;
		else obs_hash_str <= obs_hash_str;
	end



	// get the compare pin high
	always@(posedge clk) begin
		if(~resetn) cmp <= 0;
		else if(obs_hash_str==exp_hash_str) begin
			 cmp <= 1;
			 $display("XOODYAK COMPLETE!");
			 file = $fopen("output.txt","a");
			  for (k = 0; k < 32; k++) begin
				 $fwriteh(file, obs_hash_str[8*(31-k) +: 8]);
			  end
			  $fwrite(file,"\n");
			  $fclose(file);
		end
		else if (cmp) cmp <= 0;
		else cmp <= cmp;
	end
/*
initial begin
	#(150*(CLOCK_PERIOD));
	$finish();
end
*/
endmodule
