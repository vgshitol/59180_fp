`timescale 1ns / 1ps

module Testbench;

	parameter CLOCK_PERIOD = 20;
	parameter MSG_LEN = 1024;
	//parameter MSG_LEN = 19;
	
	// INPUT REGISTERS
	reg clk; 
	reg resetn; 
	reg start;
	reg load;
	reg [383:0] state_in;
	reg xoodoo_enable;
	reg [7:0] msg;
	reg [11:0] msg_len; 

	// OUTPUT REGISTERS
	wire xoodoo_complete;
	wire [383:0] state_out;
	wire [7:0] hash;
	wire [7:0] hash_len; 
	wire valid;

	// TB REGISTERS
	reg [8191:0] msg_str;
	reg [255:0] exp_hash_str;
	reg [255:0] obs_hash_str;
	reg cmp;

	reg  [255:0] test_vector [0:11] = {
		256'hEA152F2B47BCE24EFB66C479D4ADF17BD324D806E85FF75EE369EE50DC8F8BD1,
		256'h27921F8DDF392894460B70B3ED6C091E6421B7D2147DCD6031D7EFEBAD3030CC,
		256'hDD3F12E89DB41C61D3C05779705FA946A8C69C79EEFDC1B4A966A5F1AB35073D,
		256'h72ABD350DC287E8C4B95DD37BD796D79F90026C1BD4E0D99D2117BAAB26BC2CA,
		256'hA13AE46F62E433CE4CAD9E4F24C46F37B6B3815C8539A3659DAAECAAE1AB8FDB,
		256'h042383068C131A0D365B781DFCB20E855F4A68DE2072AA8D1E16181563D6F622,
		256'h415D3A751952454C1BB900700A2EB8C2814F0A30C34BC25CC37D3DE96159F4AE,
		256'h072F0834CC8FE7996E90ADED60228C18791E3A3DA38A3831DA880EDF7869909C,
		256'hC826D28C7F5BF948FBA9BB5EA028B4E377F1DE86EC5A2A1511BA4D692968EFD5,
		256'hD926F7E44B263CBA8F98E2A52B7BE175D406A2E81B462408BDBC408784C4284F,
		256'h98D44061E4D0EED4519061B947FD486B620F9B11CC3F4DF3F219E11E73B04FAD,
		256'hC23BF64CB9CE397460C685DE83EB40FE1B889CCDFDA5BE5DEA045AFCE30BB065
	};
	
	//generate clock
	always #(CLOCK_PERIOD/2) clk = ~clk;

	// Instantiate the Unit Under Test (UUT)
	XOODYAK dut1 (.clk(clk),.resetn(resetn),.start(start),.load(load),.xoodoo_complete(xoodoo_complete),.state_in(state_in),.msg(msg),
		.msg_len(msg_len),.xoodoo_enable (xoodoo_enable),.state_out(state_out),.hash(hash),.hash_len(hash_len),.valid(valid));
	
	XOODOO dut2 (.clk(clk),.resetn(resetn),.enable_xoodoo(xoodoo_enable),.state_in(state_out),.state_out(state_in),.done_permutations(xoodoo_complete));

	integer i=0,j=0,k=0;
	integer file,r;
		
	// Drive the testbench
	initial begin
		resetn=1'b1;
		clk = 1'b0;
		msg_str = 8192'h000102030405060708090A0B0C0D0E0F101112131415161718191A1B1C1D1E1F202122232425262728292A2B2C2D2E2F303132333435363738393A3B3C3D3E3F404142434445464748494A4B4C4D4E4F505152535455565758595A5B5C5D5E5F606162636465666768696A6B6C6D6E6F707172737475767778797A7B7C7D7E7F808182838485868788898A8B8C8D8E8F909192939495969798999A9B9C9D9E9FA0A1A2A3A4A5A6A7A8A9AAABACADAEAFB0B1B2B3B4B5B6B7B8B9BABBBCBDBEBFC0C1C2C3C4C5C6C7C8C9CACBCCCDCECFD0D1D2D3D4D5D6D7D8D9DADBDCDDDEDFE0E1E2E3E4E5E6E7E8E9EAEBECEDEEEFF0F1F2F3F4F5F6F7F8F9FAFBFCFDFEFF000102030405060708090A0B0C0D0E0F101112131415161718191A1B1C1D1E1F202122232425262728292A2B2C2D2E2F303132333435363738393A3B3C3D3E3F404142434445464748494A4B4C4D4E4F505152535455565758595A5B5C5D5E5F606162636465666768696A6B6C6D6E6F707172737475767778797A7B7C7D7E7F808182838485868788898A8B8C8D8E8F909192939495969798999A9B9C9D9E9FA0A1A2A3A4A5A6A7A8A9AAABACADAEAFB0B1B2B3B4B5B6B7B8B9BABBBCBDBEBFC0C1C2C3C4C5C6C7C8C9CACBCCCDCECFD0D1D2D3D4D5D6D7D8D9DADBDCDDDEDFE0E1E2E3E4E5E6E7E8E9EAEBECEDEEEFF0F1F2F3F4F5F6F7F8F9FAFBFCFDFEFF000102030405060708090A0B0C0D0E0F101112131415161718191A1B1C1D1E1F202122232425262728292A2B2C2D2E2F303132333435363738393A3B3C3D3E3F404142434445464748494A4B4C4D4E4F505152535455565758595A5B5C5D5E5F606162636465666768696A6B6C6D6E6F707172737475767778797A7B7C7D7E7F808182838485868788898A8B8C8D8E8F909192939495969798999A9B9C9D9E9FA0A1A2A3A4A5A6A7A8A9AAABACADAEAFB0B1B2B3B4B5B6B7B8B9BABBBCBDBEBFC0C1C2C3C4C5C6C7C8C9CACBCCCDCECFD0D1D2D3D4D5D6D7D8D9DADBDCDDDEDFE0E1E2E3E4E5E6E7E8E9EAEBECEDEEEFF0F1F2F3F4F5F6F7F8F9FAFBFCFDFEFF000102030405060708090A0B0C0D0E0F101112131415161718191A1B1C1D1E1F202122232425262728292A2B2C2D2E2F303132333435363738393A3B3C3D3E3F404142434445464748494A4B4C4D4E4F505152535455565758595A5B5C5D5E5F606162636465666768696A6B6C6D6E6F707172737475767778797A7B7C7D7E7F808182838485868788898A8B8C8D8E8F909192939495969798999A9B9C9D9E9FA0A1A2A3A4A5A6A7A8A9AAABACADAEAFB0B1B2B3B4B5B6B7B8B9BABBBCBDBEBFC0C1C2C3C4C5C6C7C8C9CACBCCCDCECFD0D1D2D3D4D5D6D7D8D9DADBDCDDDEDFE0E1E2E3E4E5E6E7E8E9EAEBECEDEEEFF0F1F2F3F4F5F6F7F8F9FAFBFCFDFEFF;
	    exp_hash_str = 256'hfcc4d63932d98c30cab597e60b7cca475bd9fbf984838c5cb5615c949f814615;
	   // msg_str = 8192'h000102030405060708090A0B0C0D0E0F101112;
	 	
	 	#(10*(CLOCK_PERIOD));
		resetn=1'b0;
		#(2*(CLOCK_PERIOD));
		
		resetn=1'b1;
		
		#(10*(CLOCK_PERIOD));
		for (j = 0; j < 12; j++) begin
			/* code */
			msg_len = j;
			exp_hash_str = test_vector[j];
			//#(CLOCK_PERIOD/2);
			load = 1;
			for (i=0;i<=j;i=i+1)
			begin
				msg=msg_str>>(i + 1023-j)*8;//(MSG_LEN-i-1)*8;
			//	$display("%d,%d,%x",i,j,msg);
				#(CLOCK_PERIOD);
			end
			load = 0;

			#(5*CLOCK_PERIOD);
			start = 1;
			#(CLOCK_PERIOD);
			start = 0;
			
			repeat(3000) begin
				#((CLOCK_PERIOD));
			end	
		end

		$stop;
		
	end

	// initial begin
	// 	file = $fopen("output.txt","w");
	// 	if(i) begin 
	// 		$fwrite(file,"%x\n",   hash);
	// 		i=0;
	// 	end
	// 	$fclose(file);
	// end

	
	// Get the output string
	always@(posedge clk) begin
		if(~resetn || load) obs_hash_str <= 0;
		else if(valid==1'b1) begin
		//	 $display("VALID HIGH!");
			 obs_hash_str <= {obs_hash_str[247:0],hash};
		end
		else if(obs_hash_str==exp_hash_str) obs_hash_str <= 0;
		else obs_hash_str <= obs_hash_str;
	end



	// get the compare pin high
	always@(posedge clk) begin
		if(~resetn || load) cmp <= 0;
		else if(obs_hash_str==exp_hash_str) begin
			 cmp <= 1;
			 $display("XOODYAK COMPLETE!");
			 file = $fopen("output.txt","a");
			  for (k = 0; k < 32; k++) begin
				 $fwriteh(file, obs_hash_str[8*(31-k) +: 8]);
			  end
			  $fwrite(file,"\n");
			  $fclose(file);
		end
		else if (cmp) cmp <= 0;
		else cmp <= cmp;
	end


endmodule
